// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Full Version"
// CREATED		"Fri Jun 24 17:07:43 2016"
`timescale 1ns / 1ps
`default_nettype none
  // Top level HDL module
  module maaps_daq_toplevel(
			    CK50,
			    adcfastclk_p,
			    adcframe_p,
			    spi_cs,
			    spi_sclk,
			    spi_data_in,
			    PMT_trigger,
			    adcdata_p,
			    TDC,
			    ADC_SCLK1,
			    ADC_nCS1,
			    ADCCLK1_p,
			    ADCCLK2_p,
			    L1,
			    L0,
			    spi_data_out,
			    ADC_SDIO1,
			    Z0,
			    Z0_FRAME,
			    Z0_CLK
			    );


   input wire	CK50;
   input wire	adcfastclk_p;
   input wire	adcframe_p;
   input wire	spi_cs;
   input wire	spi_sclk;
   input wire	spi_data_in;
   input wire	PMT_trigger;
   input wire [15:0] adcdata_p; // 16 serial lines
   input wire [31:0] TDC; // unused
   output wire 	     ADC_SCLK1;
   output wire 	     ADC_nCS1;
   output wire 	     ADCCLK1_p;
   output wire 	     ADCCLK2_p;
   output wire 	     L1;
   output wire 	     L0;
   output wire 	     spi_data_out;
   inout wire 	     ADC_SDIO1;
	reg rst;

   // input clock - 50 MHz 
   wire 	     sysclk;
   assign	sysclk = CK50;

   // output clocks to the two octal ADCs
   assign ADCCLK1_p = sysclk;
   assign ADCCLK2_p = sysclk;

   wire [15:0] 	     dout;
   wire 	     adc_ready; // output

   wire 	     adc_flag;
   reg [7:0] 	     adc_mode;

   // hard-wired for now
   initial adc_mode = 8'h09;
   // SPI controller to configure the external ADCs
   adc_spimaster adc_spimaster_inst(
				    .sys_clk(sysclk),
				    .reset_n(~rst),
      
				    .adc_sclk(ADC_SCLK1),
				    .adc_sdio(ADC_SDIO1),
				    .adc_cs(ADC_nCS1),
      
				    .adc_flag(adc_flag),
				    .adc_mode(adc_mode),
				    .adc_ready(adc_ready)
				    );
   
   
   
   // module to contain the input from the digitizer channels.
   // configurable how many it controls by the CHAN variable
   // howmany, offset should be made configurable - hardwired for now
   // DAVAIL and TRIGGER should also not be hardwired to their current widths.
   digi_many #(.CHAN(8)) digi_many_inst(
					.RST(rst&adc_ready), 
					.CK50(sysclk), 
					.adc_clk(adcfastclk_p), 
					.adc_frame(adcframe_p),
					.adcdata_p(adcdata_p), 
					.DOUT(dout), // output to remote
					.ZYNQ_RD_REQUEST(1),
					.howmany(8'hFF), // configuration
					.offset(8'h00), // configuration
					.DAVAIL(TDC[7:0]), // FIXME
					.TRIGGER(TDC[16:8]) // FIXME
					);

   // counter just to twiddle the LED on the digitzer
   wire [31:0] 	     dcount;
   bc_counter #(.BITS(32)) counter_inst0(
					 .CLK(sysclk),
					 .RST(rst), 
					 .BC(dcount)
					 );
   assign L0 = dcount[26]; // should be about 1 Hz
   assign L1 = dcount[25]; // should be 2x as fast as L1
   
   output wire [1:0] Z0;
   output wire 	     Z0_FRAME;
   output wire 	     Z0_CLK;

   // LVDS output to the ZYNQ
   // the Z0 clock is the slow clock; its leading edge indicates the
   // MSB of the serial output stream.
   lvds_transmitter lvds_tx_inst(
				 .DIN(dout), 
				 .CLK(sysclk),
				 .O_D(Z0),
				 .O_CLK(Z0_CLK)
				 );
   
	// self-reset on startup for now. This is a hack.
	reg [4:0] rst_cnt; 
	initial rst_cnt = 0;
	always @(posedge sysclk ) begin
		if ( rst_cnt < 31 )
			rst_cnt <= rst_cnt + 5'b1;
		if ( rst_cnt < 31) 
			rst = 1;
		else
			rst = 0;
			
	end
	
endmodule

